--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   20:10:58 04/06/2015
-- Design Name:   
-- Module Name:   C:/Users/Administrator/Desktop/xkz/TestBench.vhd
-- Project Name:  xkz
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: xkz
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TestBench IS
END TestBench;
 
ARCHITECTURE behavior OF TestBench IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT xkz_b
    PORT(
         clk : IN  std_logic;
         s5: IN std_logic;
	       s2: IN std_logic;
	       wavelength: IN std_logic_vector(8 downto 0);
         z : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal s5: std_logic := '0';
	 signal s2: std_logic := '0';
	 signal wavelength: std_logic_vector(8 downto 0) := "000000001";

 	--Outputs
   signal z : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: xkz_b PORT MAP (
          clk => clk,
          s5 => s5,
          s2 => s2,
          z => z,
          wavelength => wavelength
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- s5 process
   s5_process: process
   begin		
     s5 <= '1';
     wait for clk_period*6;
     s5 <= '0';
     wait for clk_period*1000;
   end process;
   
   
   
   -- s2 process
   s2_process: process
   begin
     wait for clk_period*6;		
     s2 <= '1';
     wait for clk_period*15;
     s2 <= '0';
     wait for clk_period*1000;
   end process;
   
   wavelength_process: process
   begin
     wait for clk_period*6;
     wait for clk_period*15;
     wavelength <= "000000001";
     wait for clk_period*10;
     wavelength <= "000000010";
     wait for clk_period*10;
     wavelength <= "000000100";
     wait for clk_period*10;
     wavelength <= "000001000";
     wait for clk_period*10;
     wavelength <= "000010000";
     wait for clk_period*10;
     wavelength <= "000100000";
     wait for clk_period*10;
     wavelength <= "001000000";
     wait for clk_period*10;
     wavelength <= "010000000";
     wait for clk_period*10;
     wavelength <= "100000000";
     wait for clk_period*9;
     wavelength <= "000000001";
     wait for clk_period*1000;
   end process;

END;
